module knight_rider();

endmodule
