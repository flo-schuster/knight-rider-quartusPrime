module knight_rider(
	input D
);



endmodule
